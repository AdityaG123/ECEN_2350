`timescale 1ns/100ps

module testbenchlab2();
reg my_ADC_CLK_10;
wire [7:0] my_HEX0, my_HEX1, my_HEX2, my_HEX3, my_HEX4, my_HEX5;
reg [1:0] my_KEY;
wire [9:0] my_LEDR;
wire [9:0] my_SW;

always
#100 my_ADC_CLK_10 = ~my_ADC_CLK_10;


toplab2test U0 (.ADC_CLK_10(my_ADC_CLK_10),.KEY(my_KEY),.SW(my_SW),.LEDR(my_LEDR),.HEX0(my_HEX0),.HEX1(my_HEX1),.HEX2(my_HEX2),.HEX3(my_HEX3),.HEX4(my_HEX4),.HEX5(my_HEX5));


initial
begin
  $dumpfile("out.vcd");
	$dumpvars;
    $display($time, " << Starting Simulation >>");
    my_ADC_CLK_10 = 0;
    my_KEY[0] = 1;
    #100000  my_KEY[0] = 0;
    #100000  my_KEY[0] = 1;
    #100000  my_KEY[0] = 0;
    #100000  my_KEY[0] = 1;
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    #100000
    $finish;
end

initial
begin
 $monitor($time,"  HEX 2: %b, HEX 1: %b, HEX 0: %b, LED: %b",my_HEX2,my_HEX1,my_HEX0,my_LEDR[1:0]);
end

endmodule
