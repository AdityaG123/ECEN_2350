module full_subtractor(Cin,a,b,diff,Cout);